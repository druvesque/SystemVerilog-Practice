class A;
    integer data;
    local integer addr;
    protected integer cmd;
    static integer cred;
endclass
