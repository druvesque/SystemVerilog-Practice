// DELTA SIMULATION TIME / CYCLE / DELAY
// SIMULATION CYCLE VS CLOCK CYCLE
// #1step, #1 <= #1step <= ##1
// 2-state variable is synthesizable?
// 

