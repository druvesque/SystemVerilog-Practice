// Verification: testing a design whether it performs the desired task and
//               measuring it's response under different stimulus.
//               Here, we focus on constrained-random, assertion based and
//               coverage-driven verification.
//               
// Testbench: piece of code that is capable of generating a wide range of
//            input test vectors for DUT and observe it's response. 
//            
//            1. Generate Stimulus
//            2. Applying Stimulus to the DUT
//            3. Capture the response
//            4. Check for correctness
//            5. Measure the progress against the overall verification goals
//            6. Convert quantity into quality
//            
// ---> SV combines the HDL and HVL features in a single language.
