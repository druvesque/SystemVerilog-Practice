// NOTES
// vlog -work work file.sv
// vsim -novopt work.tb
// vlog -help
// vsim -help
// 
// GUI
// TCL
// CORE
//
//
// Parallel Blocks in Verilog 
//
// - fork...join/join_any/join_none
// - always (always_ff, always_latch, always_comb)
// - multiple initial blocks
// - multiple parallel blocks
// - module instantiation
// - gate instantiation
// - primitive instances
// - specify blocks


