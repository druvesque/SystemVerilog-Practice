// NOTES
// vlog -work work file.sv
// vsim -novopt work.tb
// vlog -help
// vsim -help
// 
// GUI
// TCL
// CORE


