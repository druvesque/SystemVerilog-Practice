module test;

    initial begin
        $display("sizeof(int): %0d", sizeof(int));
    end
endmodule
